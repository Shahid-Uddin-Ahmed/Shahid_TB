module mux_4_to_1( 
    input [3:0] a,                 // 4-bit input called a
                       
    input [3:0] b,                 // 4-bit input called b
                       
    input [3:0] c,                 // 4-bit input called c
                       
    input [3:0] d,                 // 4-bit input called d
                       
    input [1:0] sel,               // input sel used to select between a,b,c,d
    output reg [3:0] out);         // 4-bit output based on input sel
                  
   always @ (a or b or c or d or sel) begin
      case (sel)
         2'b00 : out <= a;
         2'b01 : out <= b;
         2'b10 : out <= c;
         2'b11 : out <= d;
      endcase
   end
endmodule
